netcdf ice_shelf_v1 {
dimensions:
	ny = 40 ;
	nx = 240 ;
variables:
	double thick(ny, nx) ;
		thick:units = "m" ;
		thick:standard_name = "ice shelf thickness" ;
	double area(ny, nx) ;
		area:units = "m2" ;
		area:standard_name = "ice shelf area" ;
        double height(ny, nx) ;
                height:units = "m" ;
                height:standard_name = "location of ssh (negative if under ice shelf)" ;
}
